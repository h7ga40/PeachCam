/*
 *  TOPPERS/ASP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Advanced Standard Profile Kernel
 * 
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015,2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 * 
 *  上記著作権者は，以下の(1)～(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: tSIOPortGRPeach.cdl 1846 2019-03-28 10:22:45Z coas-nagasima $
 */

/*
 *		シリアルインタフェースドライバのターゲット依存部（GR-PEACH用）
 *		のコンポーネント記述
 */

/*
 *  GR-PEACHとRZ/A1に関する定義
 */
import_C("gr_peach.h");
import_C("device.h");

/*
 *  FIFO内蔵シリアルコミュニケーションインタフェース用 簡易SIOドライバ
 */
import("tMbedSerial.cdl");

/*
 *  シリアルインタフェースドライバのターゲット依存部の本体（シリアルイ
 *  ンタフェースドライバとSIOドライバを接続する部分）のセルタイプ
 */
celltype tSIOPortGRPeachMain {
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	[inline] entry		sSIOPort	eSIOPort;
	[optional] call		siSIOCBR	ciSIOCBR;

	/*
	 *  SIOドライバとの結合
	 */
	call			sSIOPort	cSIOPort;
	[inline] entry	siSIOCBR	eiSIOCBR;
};

/*
 *  シリアルインタフェースドライバのターゲット依存部（複合コンポーネン
 *  ト）のセルタイプ
 */
composite tSIOPortGRPeach {
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	entry				sSIOPort	eSIOPort;
	[optional] call		siSIOCBR	ciSIOCBR;

	/*
	 *  属性の定義
	 */
	attr {
		int32_t tx;								/* 送信Pin */
		int32_t rx;								/* 受信Pin */
		uint32_t	baudRate = 115200;			/* ボーレートの設定値 */
	};

	/*
	 *  SIOドライバ
	 */
	cell tMbedSerial MbedSerial {
		tx          = composite.tx;
		rx          = composite.rx;
		baudRate    = composite.baudRate;
		ciSIOCBR    = SIOPortMain.eiSIOCBR;
	};

	/*
	 *  シリアルインタフェースドライバのターゲット依存部の本体
	 */
	cell tSIOPortGRPeachMain SIOPortMain {
		ciSIOCBR            => composite.ciSIOCBR;
		cSIOPort            = MbedSerial.eSIOPort;
	};
	composite.eSIOPort => SIOPortMain.eSIOPort;
};

/*
 *  シリアルインタフェースドライバのターゲット依存部のプロトタイプ
 *
 *  サンプルプログラムが使うポートが，SIOPortTarget1に固定されているた
 *  め，ポート1とポート3を入れ換えている．具体的には，SIOPortTarget1は
 *  MbedSerialのチャネル2（チャネル番号は0から始まるので，ポート3のこと）に，
 *  SIOPortTarget3はMbedSerialのチャネル0につながっている．
 */
[prototype]
cell tSIOPortGRPeach SIOPortTarget1 {
	/* 属性の設定 */
	tx = C_EXP("P6_3");
	rx = C_EXP("P6_2");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget2 {
	/* 属性の設定 */
	tx = C_EXP("P2_5");
	rx = C_EXP("P2_6");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget3 {
	/* 属性の設定 */
	tx = C_EXP("P4_12");
	rx = C_EXP("P4_13");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget4 {
	/* 属性の設定 */
	tx = C_EXP("P2_14");
	rx = C_EXP("P2_15");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget5 {
	/* 属性の設定 */
	tx = C_EXP("P4_14");
	rx = C_EXP("P4_15");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget6 {
	/* 属性の設定 */
	tx = C_EXP("P5_3");
	rx = C_EXP("P5_4");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget7 {
	/* 属性の設定 */
	tx = C_EXP("P8_8");
	rx = C_EXP("P8_9");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget8 {
	/* 属性の設定 */
	tx = C_EXP("P5_0");
	rx = C_EXP("P5_1");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget9 {
	/* 属性の設定 */
	tx = C_EXP("P8_14");
	rx = C_EXP("P8_15");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget10 {
	/* 属性の設定 */
	tx = C_EXP("P8_13");
	rx = C_EXP("P8_11");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget11 {
	/* 属性の設定 */
	tx = C_EXP("P11_10");
	rx = C_EXP("P11_11");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget12 {
	/* 属性の設定 */
	tx = C_EXP("P6_6");
	rx = C_EXP("P6_7");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget13 {
	/* 属性の設定 */
	tx = C_EXP("P5_6");
	rx = C_EXP("P5_7");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget14 {
	/* 属性の設定 */
	tx = C_EXP("P11_1");
	rx = C_EXP("P11_2");
};

[prototype]
cell tSIOPortGRPeach SIOPortTarget15 {
	/* 属性の設定 */
	tx = C_EXP("P7_4");
	rx = C_EXP("P7_5");
};
