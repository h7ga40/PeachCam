/*
 *		C言語で記述されたアプリケーションから，TECSベースの実行時間分布
 *		集計サービスを呼び出すためのアダプタ用セルタイプの定義
 * 
 *  $Id: tHistogramAdapter.cdl 1484 2018-03-30 12:24:59Z coas-nagasima $
 */
[singleton, active]
celltype tHistogramAdapter {
	call	sHistogram		cHistogram[];
};
