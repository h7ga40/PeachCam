/*
 *		C言語で記述されたアプリケーションから，TECSベースのテストプログ
 *		ラム用サービスを呼び出すためのアダプタ用セルタイプの定義
 *
 *  $Id: tTestServiceAdapter.cdl 1428 2018-02-18 13:58:37Z coas-nagasima $
 */
[singleton, active]
celltype tTestServiceAdapter {
	call	sTestService	cTestService;
};
