/*
 *  TOPPERS/ASP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Advanced Standard Profile Kernel
 * 
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015,2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 * 
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: tSIOPortNTShell.cdl 1888 2019-04-19 09:55:29Z coas-nagasima $
 */

/*
 *		シリアルインタフェースドライバのターゲット依存部（NTShell用）
 *		のコンポーネント記述
 */

/*
 *  NTShell に関する定義
 */
import_C("termios.h");

/*
 *  SIOドライバの本体のセルタイプ
 */
celltype tSIOPortNTShellMain {
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	entry				sSIOPort		eSIOPort;
	[optional] call		siSIOCBR		ciSIOCBR;

	/*
	 *  終了処理ルーチン
	 */
	entry	sRoutineBody	eTerminate;

	attr {
		const char	*path;				/* パス名 */
	};

	var {
		bool_t			opened = false;	/* オープン済みフラグ */
		struct termios	saved_term;		/* 元の端末制御情報 */
		int_t			read_fd;		/* 読出し用ファイルディスクリプタ */
		bool_t			rcv_flag;		/* 受信文字バッファ有効フラグ */
		char			rcv_buf;		/* 受信文字バッファ */
		bool_t			rcv_rdy;		/* 受信通知コールバック許可フラグ */
		int_t			write_fd;		/* 書込み用ファイルディスクリプタ */
		bool_t			snd_flag;		/* 送信文字バッファ有効フラグ */
		char			snd_buf;		/* 送信文字バッファ */
		bool_t			snd_rdy;		/* 送信通知コールバック許可フラグ */
	};
};

/*
 *  SIOドライバ（複合コンポーネント）のセルタイプ
 */
[active]
composite tSIOPortNTShell {
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	entry				sSIOPort	eSIOPort;
	[optional] call		siSIOCBR	ciSIOCBR;

	/*
	 *  属性の定義
	 */
	attr {
		const char	*path = C_EXP("NULL");		/* パス名 */
	};

	/*
	 *  SIOドライバの本体
	 */
	cell tSIOPortNTShellMain SIOPortMain {
		path     = composite.path;
		ciSIOCBR => composite.ciSIOCBR;
	};
	composite.eSIOPort => SIOPortMain.eSIOPort;

	/*
	 *  SIOドライバの終了処理ルーチン
	 */
	cell tTerminateRoutine TerminateSIO {
		cTerminateRoutineBody = SIOPortMain.eTerminate;
	};
};
