/*
 *  TOPPERS Software
 *      Toyohashi Open Platform for Embedded Real-Time Systems
 * 
 *  Copyright (C) 2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 * 
 *  上記著作権者は，以下の(1)～(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: tHistogram.cdl 1484 2018-03-30 12:24:59Z coas-nagasima $
 */

/*
 *		実行時間分布集計サービスのコンポーネント記述ファイル
 */

import_C("syssvc/tHistogram.h");

/*
 *  実行時間分布集計サービスのシグニチャ
 */
signature sHistogram {
	/*
	 *  実行時間分布計測の初期化
   	 */
	void	initialize(void);

	/*
	 *  実行時間計測の開始
	 */
	void	beginMeasure(void);

	/*
	 *  実行時間計測の終了
	 */
	void	endMeasure(void);

	/*
	 *  実行時間分布計測の表示
	 */
	void	print(void);
};

/*
 *  実行時間分布集計サービスのセルタイプ
 */
celltype tHistogram {
	entry	sHistogram		eHistogram;

	attr {
		uint_t		maxTime = 1000;		/* 分布を記録する最大時間 */
	};
	var {
		[size_is(maxTime + 1)] uint_t	*histarea;
										/* 分布を記録するメモリ領域 */
		histtim_t	begin_time;			/* 計測開始時刻 */
		uint_t		over;				/* 最大時間を超えた度数 */
		uint_t		under;				/* 時間の逆転が疑われる度数 */
	};
};
